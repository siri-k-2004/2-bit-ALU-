module tb_alu_2bit;
 // Declare registers for inputs to the ALU (driven by test bench)
 reg [1:0] operand_a; 
 reg [1:0] operand_b; 
 reg [2:0] operation; 

 // Declare wires for outputs from the ALU (monitored by test bench)
 wire [1:0] result; 
 wire carry_out; 

 // Instantiate the 2-bit ALU module (Design Under Test - DUT)
 // Using named port connections for clarity and robustness
 alu_2bit uut(
    .operand_a(operand_a), 
    .operand_b(operand_b), 
    .operation(operation), 
    .result(result), 
    .carry_out(carry_out)
 ); 
 
 // Initial block for stimulus generation and monitoring
 initial begin
     // Enable waveform dumping for simulation tools (e.g., ModelSim)
     $dumpfile("tb_alu_2bit.vcd"); // Specify output file for waveforms
     $dumpvars(0, tb_alu_2bit); // Dump all variables in the current scope

     // Monitor inputs and outputs for changes and print to console
     $monitor("Time=%0t | OpA=%b | OpB=%b | OpCode=%b | Result=%b | CarryOut=%b", 
              $time, operand_a, operand_b, operation, result, carry_out);

     // --- Test Cases ---

     // Test Case 1: Addition (1 + 1 = 2'b10, result=00, carry=1)
     operand_a = 2'b01; 
     operand_b = 2'b01; 
     operation = 3'b000; // Addition
     #50; // Wait for 50 time units for signals to stabilize

     // Test Case 2: Subtraction (1 - 0 = 2'b01, result=01, carry=0)
     operand_a = 2'b01;
     operand_b = 2'b00;
     operation = 3'b001; // Subtraction
     #50;

     // Test Case 3: Logical AND (11 & 01 = 2'b01)
     operand_a = 2'b11; // Decimal 3
     operand_b = 2'b01; // Decimal 1
     operation = 3'b010; // Logical AND
     #50;

     // Test Case 4: Logical OR (10 | 01 = 2'b11)
     operand_a = 2'b10; // Decimal 2
     operand_b = 2'b01; // Decimal 1
     operation = 3'b011; // Logical OR
     #50;

     // Test Case 5: Logical XOR (11 ^ 10 = 2'b01)
     operand_a = 2'b11; // Decimal 3
     operand_b = 2'b10; // Decimal 2
     operation = 3'b100; // Logical XOR
     #50;

     // Test Case 6: Addition with Carry (11 + 01 = 2'b100, result=00, carry=1)
     operand_a = 2'b11; // Decimal 3
     operand_b = 2'b01; // Decimal 1
     operation = 3'b000; // Addition
     #50;

     // Test Case 7: Subtraction with Underflow (00 - 01 = 2'b11 (2's complement for -1), carry=0)
     // For unsigned operations, subtraction resulting in a negative number will wrap around.
     // The carry_out for subtraction typically indicates a borrow (0 for no borrow, 1 for borrow).
     // Here, 00 - 01 results in 11 (binary -1), and no explicit borrow flag is generated by default Verilog subtraction for unsigned.
     operand_a = 2'b00; // Decimal 0
     operand_b = 2'b01; // Decimal 1
     operation = 3'b001; // Subtraction
     #50;

     // Test Case 8: All zeros for logical operations (00 & 00 = 00, 00 | 00 = 00, 00 ^ 00 = 00)
     operand_a = 2'b00;
     operand_b = 2'b00;
     operation = 3'b010; // AND
     #50;
     operation = 3'b011; // OR
     #50;
     operation = 3'b100; // XOR
     #50;

     // Test Case 9: Max values for logical operations (11 & 11 = 11, 11 | 11 = 11, 11 ^ 11 = 00)
     operand_a = 2'b11;
     operand_b = 2'b11;
     operation = 3'b010; // AND
     #50;
     operation = 3'b011; // OR
     #50;
     operation = 3'b100; // XOR
     #50;

     // End simulation
     #100 $finish; 
 end
endmodule
